
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h81868106,
    32'h82868206,
    32'h83868306,
    32'h84868406,
    32'h85868506,
    32'h86868606,
    32'h87868706,
    32'h88868806,
    32'h89868906,
    32'h8A868A06,
    32'h8B868B06,
    32'h8C868C06,
    32'h8D868D06,
    32'h8E868E06,
    32'h8F868F06,
    32'h000FC117,
    32'hF3010113,
    32'h00000D17,
    32'h470D0D13,
    32'h00000D97,
    32'h468D8D93,
    32'h01BD5763,
    32'h000D2023,
    32'hDDE30D11,
    32'h0513FFAD,
    32'h05930000,
    32'h00EF0000,
    32'h00003080,
    32'h00A5C7B3,
    32'h0037F793,
    32'h00C50733,
    32'h00079663,
    32'h00300793,
    32'h02C7E463,
    32'h00050793,
    32'h00E56C63,
    32'h00008067,
    32'h0005C683,
    32'h00178793,
    32'h00158593,
    32'hFED78FA3,
    32'hFEE7E8E3,
    32'h00008067,
    32'h00357793,
    32'h08079263,
    32'h00050793,
    32'hFFC77693,
    32'hFE068613,
    32'h08C7F663,
    32'h0005A383,
    32'h0045A283,
    32'h0085AF83,
    32'h00C5AF03,
    32'h0105AE83,
    32'h0145AE03,
    32'h0185A303,
    32'h01C5A883,
    32'h02458593,
    32'h02478793,
    32'hFFC5A803,
    32'hFC77AE23,
    32'hFE57A023,
    32'hFFF7A223,
    32'hFFE7A423,
    32'hFFD7A623,
    32'hFFC7A823,
    32'hFE67AA23,
    32'hFF17AC23,
    32'hFF07AE23,
    32'hFADFF06F,
    32'h0005C683,
    32'h00178793,
    32'h00158593,
    32'hFED78FA3,
    32'h0037F693,
    32'hFE0696E3,
    32'hF89FF06F,
    32'h00050793,
    32'hFF1FF06F,
    32'h0005A603,
    32'h00478793,
    32'h00458593,
    32'hFEC7AE23,
    32'hFED7E8E3,
    32'hF4E7EAE3,
    32'h00008067,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h66211141,
    32'h001105B7,
    32'hC6064501,
    32'h87B73DF5,
    32'h07370011,
    32'hB6B70010,
    32'hA8030011,
    32'h43C80007,
    32'h47D0478C,
    32'h01072023,
    32'hC70CC348,
    32'h07C1C750,
    32'h94E30741,
    32'h77B7FED7,
    32'hA4231A10,
    32'h07930007,
    32'h80670800,
    32'h00010007,
    32'h00010001,
    32'h450140B2,
    32'h80820141,
    32'h1B0057B7,
    32'h11014798,
    32'hCE0676C1,
    32'hCA26CC22,
    32'hC64EC84A,
    32'hC256C452,
    32'h8F75C05A,
    32'h4BD8C798,
    32'h000706B7,
    32'hFFF80637,
    32'hCBD88F55,
    32'h06B74FD8,
    32'h16FDFFF9,
    32'hCFD88F75,
    32'h06B74FD8,
    32'h167D0008,
    32'hCFD88F55,
    32'h46814BD8,
    32'h8F7145A1,
    32'hC7B7CBD8,
    32'h47111A12,
    32'hC3D84601,
    32'h0FF00513,
    32'h458122E9,
    32'h22ED4501,
    32'h2ADD4501,
    32'h45054581,
    32'h24316441,
    32'h4485147D,
    32'h8D612425,
    32'hFE951EE3,
    32'h46014681,
    32'h451145A1,
    32'h4581224D,
    32'h22C94501,
    32'h22F94501,
    32'h45054581,
    32'h22D56441,
    32'h4485147D,
    32'h8D612401,
    32'hFE951EE3,
    32'hFF0104B7,
    32'h00FF0437,
    32'h69854901,
    32'hF0048493,
    32'h0FF40413,
    32'h161346E1,
    32'h45A10089,
    32'h2295450D,
    32'h45014581,
    32'h65212251,
    32'h45812A41,
    32'h22654501,
    32'h854A65A1,
    32'h86CA2AD1,
    32'h01390633,
    32'h06914298,
    32'h00871793,
    32'h8F618321,
    32'h8FD98FE5,
    32'h01079713,
    32'h8FD983C1,
    32'hFEF6AE23,
    32'hFED612E3,
    32'h67A1994E,
    32'hFAF91AE3,
    32'h147D6441,
    32'h22794485,
    32'h1EE38D61,
    32'h09B7FE95,
    32'h0937FF01,
    32'h0AB700FF,
    32'h0A370080,
    32'h6B050010,
    32'hF0098993,
    32'h0FF90913,
    32'h001004B7,
    32'h00103437,
    32'h865646E1,
    32'h450D45A1,
    32'h458120DD,
    32'h22194501,
    32'h2A096521,
    32'h45014581,
    32'h65A1222D,
    32'h2A998552,
    32'h063386D2,
    32'h4298016A,
    32'h17930691,
    32'h83210087,
    32'h01277733,
    32'h0137F7B3,
    32'h97138FD9,
    32'h83C10107,
    32'hAE238FD9,
    32'h90E3FEF6,
    32'h9A5AFEC6,
    32'h19E39AA6,
    32'h77B7FA8A,
    32'hA4231A10,
    32'h07930007,
    32'h80670800,
    32'h00010007,
    32'h00010001,
    32'h446240F2,
    32'h494244D2,
    32'h4A2249B2,
    32'h4B024A92,
    32'h61054501,
    32'h67C18082,
    32'h17FD1101,
    32'hC63ECE06,
    32'h17FD47B2,
    32'hFFEDC63E,
    32'h1A1077B7,
    32'hCB8947DC,
    32'h89634705,
    32'h352D00E7,
    32'h450140F2,
    32'h80826105,
    32'hBFDD33F1,
    32'h001187B7,
    32'h00100737,
    32'h0011B6B7,
    32'h0007A803,
    32'h478C43C8,
    32'h202347D0,
    32'hC3480107,
    32'hC750C70C,
    32'h074107C1,
    32'hFED794E3,
    32'h001107B7,
    32'h1A107737,
    32'h8793C71C,
    32'h80670807,
    32'h00010007,
    32'h00010001,
    32'h0793BF55,
    32'h8F8D0200,
    32'h00F51533,
    32'hC7376791,
    32'h06A21A12,
    32'hF0078793,
    32'h8EFDC708,
    32'h03F5F593,
    32'h8ECDC750,
    32'h8082CB14,
    32'h05C20542,
    32'h8DC98141,
    32'h1A12C7B7,
    32'h8082CBCC,
    32'h1A12C737,
    32'h11414B1C,
    32'hC63E0542,
    32'h07C247B2,
    32'h8D5D83C1,
    32'h47B2C62A,
    32'h0141CB1C,
    32'h47858082,
    32'h95B305A1,
    32'h953300B7,
    32'h678500A7,
    32'hF0078793,
    32'h75138DFD,
    32'h8DC90FF5,
    32'h1A12C7B7,
    32'h8082C38C,
    32'h1A12C7B7,
    32'h1141439C,
    32'h4532C63E,
    32'h80820141,
    32'h4055D793,
    32'hF7931141,
    32'hC43E7FF7,
    32'hC58189FD,
    32'h078547A2,
    32'hC602C43E,
    32'h47A24732,
    32'h02F75563,
    32'h1A12C737,
    32'h87C1431C,
    32'h0FF7F793,
    32'h47B2DFE5,
    32'h46B2530C,
    32'h97AA078A,
    32'hC6360685,
    32'h46A24632,
    32'h41E3C38C,
    32'h0141FED6,
    32'h00008082,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule