    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    00000013
    0100006F
    0100006F
    0080006F
    0040006F
    0000006F
    00000093
    81868106
    82868206
    83868306
    84868406
    85868506
    86868606
    87868706
    88868806
    89868906
    8A868A06
    8B868B06
    8C868C06
    8D868D06
    8E868E06
    8F868F06
    000FC117
    F3010113
    00000D17
    46CD0D13
    00000D97
    464D8D93
    01BD5763
    000D2023
    DDE30D11
    0513FFAD
    05930000
    00EF0000
    00003060
    00A5C7B3
    0037F793
    00C50733
    00079663
    00300793
    02C7E463
    00050793
    00E56C63
    00008067
    0005C683
    00178793
    00158593
    FED78FA3
    FEE7E8E3
    00008067
    00357793
    08079263
    00050793
    FFC77693
    FE068613
    08C7F663
    0005A383
    0045A283
    0085AF83
    00C5AF03
    0105AE83
    0145AE03
    0185A303
    01C5A883
    02458593
    02478793
    FFC5A803
    FC77AE23
    FE57A023
    FFF7A223
    FFE7A423
    FFD7A623
    FFC7A823
    FE67AA23
    FF17AC23
    FF07AE23
    FADFF06F
    0005C683
    00178793
    00158593
    FED78FA3
    0037F693
    FE0696E3
    F89FF06F
    00050793
    FF1FF06F
    0005A603
    00478793
    00458593
    FEC7AE23
    FED7E8E3
    F4E7EAE3
    00008067
    00000000
    00000000
    00000000
    00000000
    66211141
    001105B7
    C6064501
    87B73DF5
    07370011
    B6B70010
    A8030011
    43C80007
    47D0478C
    01072023
    C70CC348
    07C1C750
    94E30741
    77B7FED7
    A4231A10
    07930007
    80670800
    00010007
    00010001
    450140B2
    80820141
    1B0057B7
    11014798
    CE0676C1
    CA26CC22
    C64EC84A
    C256C452
    8F75C05A
    4BD8C798
    000706B7
    FFF80637
    CBD88F55
    06B74FD8
    16FDFFF9
    CFD88F75
    06B74FD8
    167D0008
    CFD88F55
    46814BD8
    8F7145A1
    C7B7CBD8
    47111A12
    C3D84601
    0FF00513
    458122E1
    22E54501
    2AD54501
    45054581
    24296441
    4485147D
    8D61241D
    FE951EE3
    46014681
    451145A1
    45812245
    22C14501
    22F14501
    45054581
    22CD6441
    4485147D
    8D612AFD
    FE951EE3
    FF0104B7
    00FF0437
    69854901
    F0048493
    0FF40413
    161346E1
    45A10089
    228D450D
    45014581
    65212249
    45812279
    225D4501
    854A65A1
    86CA2AC9
    01390633
    06914298
    00871793
    8F618321
    8FD98FE5
    01079713
    8FD983C1
    FEF6AE23
    FED612E3
    67A1994E
    FAF91AE3
    147D6441
    22714485
    1EE38D61
    09B7FE95
    0937FF01
    0AB700FF
    0A370080
    6B050010
    F0098993
    0FF90913
    001004B7
    00103437
    865646E1
    450D45A1
    458120D5
    22114501
    2A016521
    45014581
    65A12225
    2A918552
    063386D2
    4298016A
    17930691
    83210087
    01277733
    0137F7B3
    97138FD9
    83C10107
    AE238FD9
    90E3FEF6
    9A5AFEC6
    19E39AA6
    77B7FA8A
    A4231A10
    07930007
    80670800
    00010007
    00010001
    446240F2
    494244D2
    4A2249B2
    4B024A92
    80826105
    110167C1
    CE0617FD
    47B2C63E
    C63E17FD
    77B7FFED
    47DC1A10
    4705CB89
    00E78963
    40F23535
    61054501
    33F98082
    87B7BFDD
    07370011
    B6B70010
    A8030011
    43C80007
    47D0478C
    01072023
    C70CC348
    07C1C750
    94E30741
    07B7FED7
    77370011
    C71C1A10
    08078793
    00078067
    00010001
    BF550001
    02000793
    15338F8D
    679100F5
    1A12C737
    879306A2
    C708F007
    F5938EFD
    C75003F5
    CB148ECD
    05428082
    814105C2
    C7B78DC9
    CBCC1A12
    C7378082
    4B1C1A12
    05421141
    47B2C63E
    83C107C2
    C62A8D5D
    CB1C47B2
    80820141
    05A14785
    00B795B3
    00A79533
    87936785
    8DFDF007
    0FF57513
    C7B78DC9
    C38C1A12
    C7B78082
    439C1A12
    C63E1141
    01414532
    D7938082
    11414055
    7FF7F793
    89FDC43E
    47A2C581
    C43E0785
    4732C602
    556347A2
    C73702F7
    431C1A12
    F79387C1
    DFE50FF7
    530C47B2
    078A46B2
    068597AA
    4632C636
    C38C46A2
    FED641E3
    80820141
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
    00000000
