`define USE_VLOG
// `define MEM_INIT_ZERO
// `define SIMULATION



